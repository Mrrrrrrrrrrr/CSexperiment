`include "lib/defines.vh"
module CTRL(
    input wire rst,
    input wire stallreq_for_ex,
    input wire stallreq_for_load,

    // output reg flush,
    // output reg [31:0] new_pc,
    output reg [`StallBus-1:0] stall
);  
    always @ (*) begin
        if (rst) begin
            stall = `StallBus'b0;
        end
        else begin
            stall = stallreq_for_load ? `StallBus'b000111 :
                    stallreq_for_ex ? `StallBus'b001111 :
                    `StallBus'b0;
        end
    end

endmodule